`timescale 1ns / 1ps // �������ʱ�䵥λΪ1ns������Ϊ1ps
module tb_TBS_TX;
    // -- �������� --
    localparam CLK_FREQ    = 50_000_000;
    localparam BAUD_RATE   = 115200;
    localparam CLK_PERIOD  = 1_000_000_000 / CLK_FREQ; // 20ns
    localparam BIT_PERIOD  = 1_000_000_000 / BAUD_RATE; // ~8680ns
    // -- �źŶ��� --
    reg clk_50M;
    reg rst_n;
    reg rs232_in; // DUT ����
    wire TBS_out;  // DUT ���
    
    //----------------------------------------------------------------
    // ��������ģ�� (DUT)
    //----------------------------------------------------------------
    TBS_TX #(
        .CLK_FREQ(CLK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) u_tbs_tx (
        .clk_50M(clk_50M),
        .rst_n(rst_n),
        .rs232_in(rs232_in),
        .TBS_out(TBS_out)
    );
    //----------------------------------------------------------------
    // 1. ʱ�Ӻ͸�λ��������
    //----------------------------------------------------------------
    // ����ʱ��
    initial begin
        clk_50M = 0;
        forever #(CLK_PERIOD / 2) clk_50M = ~clk_50M;
    end
    // ���ɸ�λ�źźͲ���������
    initial begin
        // ��ʼ���͸�λ
        rst_n = 1'b0;
        rs232_in = 1'b1; // RS-232 ����Ϊ��
        #200;
        rst_n = 1'b1;
        #200;
        $display("------------------- Simulation Start -------------------");
        
        // �������񣬷��Ͳ�������
        send_rs232_byte(8'h55); // ���� 01010101
        send_rs232_byte(8'hA3); // ���� 10100011
        send_rs232_byte(8'h01); // ���� 00000001
        send_rs232_byte(8'h06); // ���� 00000110
        send_rs232_byte(8'h0B); // ���� 00001100
        send_rs232_byte(8'h0F); // ���� 00001111
        send_rs232_byte(8'h6B); // ���� 01101100
        send_rs232_byte(8'hBB); // ���� 11001100
        send_rs232_byte(8'hFB); // ���� 11111100
        send_rs232_byte(8'h00); // ����ȫ 0
        send_rs232_byte(8'hFF); // ����ȫ 1
        
        #1_000_000;
        
        $display("------------------- Simulation Finish -------------------");
        $finish;
    end
    //----------------------------------------------------------------
    // 2. ������������ (Stimulus)
    //----------------------------------------------------------------
    // ����һ���������ڷ���һ���ֽڵı�׼ RS-232 ��ʽ����
    task send_rs232_byte;
        input [7:0] data_to_send;
        integer i;
        begin
            $display("At time %0t ns, sending RS232 byte: 0x%h", $time, data_to_send);
            
            // -- ������ʼλ (�͵�ƽ������һ����������) --
            rs232_in = 1'b0;
            #(BIT_PERIOD);
            // -- ����8λ����λ (�ӵ�λ����λ) --
            for (i = 0; i < 8; i = i + 1) begin
                rs232_in = data_to_send[i];
                #(BIT_PERIOD);
            end
            // -- ����ֹͣλ (�ߵ�ƽ������һ����������) --
            rs232_in = 1'b1;
            #(BIT_PERIOD);
            
            // �����ֽ�֮������һЩ����ʱ��
            #(BIT_PERIOD * 20);
        end
    endtask
    //----------------------------------------------------------------
    // 3. ��غͱȽ� (Monitor)
    //----------------------------------------------------------------
    // ��عؼ��ź�
    initial begin
        $monitor("At time %0t ns: rst_n=%b, rs232_in=%b ===> TBS_out=%b",
                 $time, rst_n, rs232_in, TBS_out);
    end
endmodule
    