module ortho_square
#(
    parameter FREQ_DIV = 250_000      // �����ڼ���ֵ�����ⲿ����ʱ����
)
(
    input  wire clk_50M,             // ϵͳʱ��
    input  wire rst_n,           // �͵�ƽ�첽��λ
    output reg  sq_0deg,         // 0�� ����
    output reg  sq_90deg         // 90�� ����
);

// ������λ���Զ�����
localparam CTR_WIDTH = $clog2(FREQ_DIV);
reg [CTR_WIDTH-1:0] cnt;

// �������߼�
always @(posedge clk_50M or negedge rst_n) begin
    if (!rst_n) begin
        cnt <= 0;
    end
    else if (cnt == FREQ_DIV - 1) begin
        cnt <= 0;
    end
    else begin
        cnt <= cnt + 1'b1;
    end
end

// 0�� �����������ڷ�ת
always @(posedge clk_50M or negedge rst_n) begin
    if (!rst_n)
        sq_0deg <= 1'b0;
    else if (cnt == FREQ_DIV - 1)
        sq_0deg <= ~sq_0deg;
end


always @(posedge clk_50M or negedge rst_n) begin
    if (!rst_n)
        sq_90deg <= 1'b0;
    else if (cnt == (FREQ_DIV >> 1) - 1)
        sq_90deg <= ~sq_90deg;
end

endmodule
