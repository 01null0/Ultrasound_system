`timescale 1ns / 1ps

module tb_UART_TX();
    // �����ź�
    reg clk_50M;
    reg rst_n;
    reg [11:0] ad_data;
    reg ad_done;
    
    // ����ź�
    wire rs232_tx;

    wire [5:0]test_bit_cnt;
    
    // ʵ����UART_TXģ��
    UART_TX uut (
        .clk_50M(clk_50M),
        .rst_n(rst_n),
        .ad_data(ad_data),
        .ad_done(ad_done),

        
        .test_bit_cnt(test_bit_cnt),

        .rs232_tx(rs232_tx)
    );
    
    // ʱ�����ɣ�50MHz
    always #10 clk_50M = ~clk_50M;
    
    // ��������
    initial begin
        // ��ʼ���ź�
        clk_50M = 0;
        rst_n = 0;
        ad_data = 12'h000;
        ad_done = 0;
        
        // ��λ
        #100 rst_n = 1;
        
        // ����1����������
        #100 ad_data = 12'hABC;
        ad_done = 1;
        #20 ad_done = 0;
        
        // �ȴ��������
        #1_000_000; // �ȴ��㹻��ʱ����ȷ���������
        
        // ����2��������һ������
        #100 ad_data = 12'h123;
        ad_done = 1;
        #20 ad_done = 0;
        
        // �ȴ��������
        #1_000_000;

        // ����3��������һ������
        #100 ad_data = 12'h001;
        ad_done = 1;
        #20 ad_done = 0;
        
        // �ȴ��������
        #1_000_000;
        // ����4��������һ������
        #100 ad_data = 12'h017;
        ad_done = 1;
        #20 ad_done = 0;
        
        // �ȴ��������
        #1_000_000;
        
        // ��������
        #100 $finish;
    end
    
    // ������
    initial begin
        $monitor("Time = %t, TX = %b, ad_data = %h, ad_done = %b", 
                 $time, rs232_tx, ad_data, ad_done);
    end
endmodule