module TBS_TX #(
    // -- ���������� --
    parameter CLK_FREQ    = 50_000_000, // ϵͳʱ��Ƶ�� (��λ: Hz)
    parameter BAUD_RATE   = 115200      // �����Ĳ�����
) (
    input                       clk_50M,        // ϵͳʱ��
    input                       rst_n,      // �첽��λ���͵�ƽ��Ч

    // -- ��׼ UART �ӿ� --
    input                       rs232_in,   // ���Ա�׼ UART_TX ģ�������ź�

    // -- TBS ���߽ӿ� --
    output                      TBS_out     // ����� TBS ����
);

    // UART_TX/RX �� BAUD_CNT_MAX = 434����ʾ 435 ��ʱ�����ڡ�
    localparam BIT_PERIOD_COUNT  = 434; // �޸���Ӳ����Ϊ 434����ʹ�� (CLK_FREQ / BAUD_RATE) + 1 ����ȷ�������߼�

    localparam PULSE_WIDTH_COUNT = BIT_PERIOD_COUNT / 10; // �����ȶ���Ϊ�������ڵ� 10%
    // ��ȷλ����㣬$clog2(N) - 1 ��ָ N ��ֵ (0��N-1) ��������λ����
    localparam PULSE_CNT_WIDTH   = $clog2(PULSE_WIDTH_COUNT) - 1;
    localparam BAUD_CNT_WIDTH    = $clog2(BIT_PERIOD_COUNT) - 1;
    
    //----------------------------------------------------------------
    // �ڲ��źŶ���
    //----------------------------------------------------------------
    // -- ����������� --
    reg [PULSE_CNT_WIDTH:0] pulse_cnt;  

    // -- ����ͬ������ؼ�� --
    reg                 rs232_in_sync_d1;
    reg                 rs232_in_sync_d2;
    wire                start_of_frame_detected; // ֡��ʼ�½��ؼ��

    // -- ������ʱ�Ӻ�״̬���� --
    reg [BAUD_CNT_WIDTH:0]  baud_cnt;         
    reg [3:0]               bit_cnt;         // ����λ������ (0-9, ��Ӧ��ʼλ, 8*����λ, ֹͣλ)
    reg                     tx_active;       // ֡���伤��״̬��־
    wire                    baud_tick;       // ���������壬��־��һ���������ڵĽ���
    
    // ����10�����ӳٵ���λ�Ĵ���
    reg [9:0]               baud_tick_delay_sr; 

    //----------------------------------------------------------------
    // �����ź�ͬ�� �� ���ؼ��
    //----------------------------------------------------------------
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            rs232_in_sync_d1 <= 1'b1;
            rs232_in_sync_d2 <= 1'b1;
        end else begin
            rs232_in_sync_d1 <= rs232_in;
            rs232_in_sync_d2 <= rs232_in_sync_d1;
        end
    end

    // ���� tx δ����ʱ���½��زű���Ϊ��֡�Ŀ�ʼ
    assign start_of_frame_detected = rs232_in_sync_d2 & ~rs232_in_sync_d1 & ~tx_active;
    
    //----------------------------------------------------------------
    // �����ʽ�������״̬��
    //----------------------------------------------------------------
    // �����ʼ�����
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            baud_cnt <= 0;
        end else if (tx_active) begin
            if (baud_cnt == BIT_PERIOD_COUNT - 1) begin
                baud_cnt <= 0;
            end else begin
                baud_cnt <= baud_cnt + 1;
            end
        end else begin
            baud_cnt <= 0;
        end
    end
    
    // ��ÿ���������ڵı߽����һ�������ڵ� tick �ź�
    assign baud_tick = (tx_active && (baud_cnt == BIT_PERIOD_COUNT - 1));

    // ����״̬��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            tx_active <= 1'b0;
            bit_cnt   <= 0;
        end else begin
            if (start_of_frame_detected) begin
                tx_active <= 1'b1;
                bit_cnt   <= 0; // ׼����ʼ��������ʼλ�ǵ�0����
            end else if (baud_tick) begin
                if (bit_cnt == 9) begin // ����1λֹͣλ����10��bit (0-9)
                    tx_active <= 1'b0;
                    bit_cnt   <= 0;
                end else begin
                    bit_cnt <= bit_cnt + 1;
                end
            end
        end
    end
    
    //----------------------------------------------------------------
    // 10�����ӳٲ������Ա���ʱ����
    // baud_tick ������ǰһ���������ڵĽ�����
    // baud_tick_d10 ���ڵ�ǰ�������ڵĿ�ʼ�� 10 ��ʱ�������ڷ�����
    // �ṩһ���ȶ��Ĳ����㡣
    //----------------------------------------------------------------
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            baud_tick_delay_sr <= 10'b0;
        end else begin
            // �� baud_tick ������λ�Ĵ��������λ�����������λ�ƶ�
            baud_tick_delay_sr <= {baud_tick_delay_sr[8:0], baud_tick};
        end
    end

    // �����ӳ�10�ĺ���źţ�ȡ��λ�Ĵ��������λ
    wire baud_tick_d10 = baud_tick_delay_sr[9];

    //----------------------------------------------------------------
    // �������ɴ����߼�
    //----------------------------------------------------------------
    // ���崥��������
    // 1. ֡�Ŀ�ʼ (start_of_frame_detected) - ����ʼλ������Ӧ��
    // 2. �ڱ������ڱ߽��10�� (baud_tick_d10)�����Ҵ�ʱ����������Ϊ�͵�ƽ - ȷ������λ�������ȶ��ԡ�
    // ���ֻ�ϴ����Ǻ���ģ���ʼλ�½���������ȷ��֡��ʼ�źţ�Ӧ������Ӧ��
    // ����������λ����Ҫ���ȶ��Ĳ����㡣
    wire trigger_pulse = start_of_frame_detected ||
                         (tx_active && baud_tick_d10 && (rs232_in_sync_d1 == 1'b0)); // ������baud_tick_d10ֻ��tx_activeʱ�Ų���

    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            pulse_cnt <= PULSE_WIDTH_COUNT;
        end else if (trigger_pulse) begin
            pulse_cnt <= 0;
        end else if (pulse_cnt < PULSE_WIDTH_COUNT) begin
            pulse_cnt <= pulse_cnt + 1'b1;
        end else begin
            pulse_cnt <= PULSE_WIDTH_COUNT;
        end
    end
    
    //----------------------------------------------------------------
    // ����ź����� (�˲����߼�����)
    //----------------------------------------------------------------
    assign TBS_out = (pulse_cnt < PULSE_WIDTH_COUNT) ? 1'b0 : 1'b1;

endmodule
