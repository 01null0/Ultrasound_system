module TBS_RX #(
    // -- ���������� --
    parameter CLK_FREQ    = 50_000_000, // ϵͳʱ��Ƶ�� (��λ: Hz)
    parameter BAUD_RATE   = 115200      // �����Ĳ�����
) (
    input                       clk_50M,        // ϵͳʱ��
    input                       rst_n,      // �첽��λ���͵�ƽ��Ч

    // -- TBS ���߽ӿ� --
    input                       TBS_in,     // ���� TBS ���ߵ������ź�

    // -- ��׼ UART �ӿ� --
    output                      rs232_out   // �������׼ UART_RX ģ��������
);

    //----------------------------------------------------------------
    // ���ز�������
    //----------------------------------------------------------------
    // ����ÿ���������ڶ�Ӧ��ʱ����������
    // localparam BIT_PERIOD_COUNT = CLK_FREQ / BAUD_RATE;
    localparam BIT_PERIOD_COUNT = 434;
    // Ϊ���������������λ��ʹ�� $clog2 ���Ż���Դ��45
    localparam CNT_WIDTH = $clog2(BIT_PERIOD_COUNT);

    //----------------------------------------------------------------
    // �ڲ��źŶ���
    //----------------------------------------------------------------
    reg  [CNT_WIDTH:0]  stretch_cnt;        // ������������ļ�����
    reg                 tbs_in_sync_d1;     // ����ͬ���Ĵ�������һ��
    reg                 tbs_in_sync_d2;     // ����ͬ���Ĵ������ڶ���
    wire                falling_edge_detected; // �½��ؼ���־

    //----------------------------------------------------------------
    // �����ź�ͬ�� �� ���ؼ��
    //----------------------------------------------------------------
    // ���첽�� TBS_in �����ź�ͬ����ϵͳʱ�����Է�ֹ����̬���⡣
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            tbs_in_sync_d1 <= 1'b1;
            tbs_in_sync_d2 <= 1'b1;
        end else begin
            tbs_in_sync_d1 <= TBS_in;
            tbs_in_sync_d2 <= tbs_in_sync_d1;
        end
    end

    // ��ͬ������ź��ϼ���½��ء��½��ر�־��һ�� '0' ���صĿ�ʼ��
    assign falling_edge_detected = tbs_in_sync_d2 & ~tbs_in_sync_d1;

    //----------------------------------------------------------------
    // ������������߼�
    //----------------------------------------------------------------
    // ����⵽�½���ʱ���˼����������㲢��ʼΪһ�������ı������ڼ�ʱ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            stretch_cnt <= BIT_PERIOD_COUNT;
        end else if (falling_edge_detected) begin
            // һ�� '0' ���ص�����������ʱ������ʼ���졣
            stretch_cnt <= 0;
        end else if (stretch_cnt < BIT_PERIOD_COUNT) begin
            // ��һ�����������ڳ���������
            stretch_cnt <= stretch_cnt + 1'b1;
        end else begin
            // ����״̬���ʱ�����󣬽�������������ֵ���ȴ���һ�δ�����
            stretch_cnt <= BIT_PERIOD_COUNT;
        end
    end

    //----------------------------------------------------------------
    // ����ź�����
    //----------------------------------------------------------------
    // ֻҪ����������ڹ��� (����ֵС�ڱ�������)������ͱ���Ϊ�͵�ƽ��
    // �������Ϊ�ߵ�ƽ (����״̬)��
    assign rs232_out = (stretch_cnt < BIT_PERIOD_COUNT) ? 1'b0 : 1'b1;

endmodule
