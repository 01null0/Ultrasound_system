`timescale 1ns / 1ps

module tb_Ultrasound_system;

    // ============================================================
    // 1. �źŶ���
    // ============================================================
    reg  clk_50M;
    reg  rst_n;
    reg  TBS_in;  // ���룺TBS Э������
    reg  ad_in;  // ���룺ģ�� AD7352 �Ĵ���������� (SDATA)

    // ����ź�
    wire TBS_out;
    wire ad_cs;
    wire ad_clk;
    wire relay;
    wire VIN_1, VIN_2, VIN_3, VIN_4;

    // ============================================================
    // 2. ��������
    // ============================================================
    parameter CLK_FREQ = 50_000_000;
    parameter BAUD_RATE = 115200;
    parameter BIT_PERIOD = 1000000000 / BAUD_RATE;  // ~8680ns
    parameter PULSE_WIDTH = BIT_PERIOD / 8;  // TBS խ������

    // ============================================================
    // 3. ʵ��������ģ��
    // ============================================================
    Ultrasound_system u_dut (
        .clk_50M(clk_50M),
        .rst_n  (rst_n),
        .TBS_in (TBS_in),
        .ad_in  (ad_in),
        .TBS_out(TBS_out),
        .ad_cs  (ad_cs),
        .ad_clk (ad_clk),
        .relay  (relay),
        .VIN_1  (VIN_1),
        .VIN_2  (VIN_2),
        .VIN_3  (VIN_3),
        .VIN_4  (VIN_4)
    );

    // ============================================================
    // 4. ���ؼ��������ض��� Order_4s �����Լ��ٷ���
    //    ���뼶/���뼶������С���Ա��ڶ�ʱ���ڹ۲쵽������ AD �ɼ�����
    // ============================================================
    // 4�� -> ��Ϊ 1ms (�㹻������)
    // defparam u_dut.inst4_Order_4s.Time_4s = 32'd50_000;

    // // 10ms -> ��Ϊ 200us (10000��ʱ��)�����̳�ʼ�ȴ�ʱ��
    // defparam u_dut.inst4_Order_4s.Time_10ms = 19'd10_000;

    // // 6ms -> ��Ϊ 100us (5000��ʱ��)��AD �������ڳ���
    // defparam u_dut.inst4_Order_4s.Time_6ms = 19'd5_000;

    // // 3ms -> ��Ϊ 50us (2500��ʱ��)������ä���ȴ�ʱ��
    // defparam u_dut.inst4_Order_4s.Time_3ms = 19'd2_500;

    // // 1us -> ��Ϊ 50��ʱ�� (���� 1MHz �����ʲ��䣬��֤ SPI ʱ����ȷ)
    // defparam u_dut.inst4_Order_4s.Time_1us = 16'd50;

    // ============================================================
    // 5. �ź�̽�� (Debug Signals)
    // ============================================================
    wire [ 2:0] debug_command = u_dut.inst3_UART_RX.command;
    wire [ 2:0] debug_uart_state = u_dut.inst3_UART_RX.state;
    //Order_4S ״̬
    wire        debug_Exc_start = u_dut.inst4_Order_4s.Exc_start;
    wire [ 2:0] debug_current_state = u_dut.inst4_Order_4s.current_state;
    // �۲� AD ������������
    wire [11:0] debug_ad_out_data = u_dut.inst9_AD.ad_out;
    wire        debug_ad_done = u_dut.inst9_AD.ad_done;
    //���������
    wire [11:0] debug_fifo_q = u_dut.inst_Echo_Correlation.fifo_q;
    wire [19:0] debug_echo_tof = u_dut.inst_Echo_Correlation.echo_tof;

    //wire debug_c0=u_dut.inst6_pll.c0;

    // ============================================================
    // 6. ʱ������
    // ============================================================
    initial begin
        clk_50M = 0;
        forever #10 clk_50M = ~clk_50M;  // 20ns ���� (50MHz)
    end

    // ============================================================
    // 7. ���񣺷��� TBS ����
    // ============================================================
    task send_tbs_byte;
        input [7:0] data;
        integer k;
        begin
            // Start Bit (Low Pulse)
            TBS_in = 0;
            #(PULSE_WIDTH);
            TBS_in = 1;
            #(BIT_PERIOD - PULSE_WIDTH);
            // Data Bits (LSB First)
            for (k = 0; k < 8; k = k + 1) begin
                if (data[k] == 1'b0) begin
                    TBS_in = 0;
                    #(PULSE_WIDTH);
                    TBS_in = 1;
                    #(BIT_PERIOD - PULSE_WIDTH);
                end
                else begin
                    TBS_in = 1;
                    #(BIT_PERIOD);
                end
            end
            // Stop Bit
            TBS_in = 1;
            #(BIT_PERIOD);
            // Inter-frame gap
            #(BIT_PERIOD * 2);
        end
    endtask

    // ============================================================
    // 8. AD7352 ��Ϊģ�� (��ȡ ad_data.hex ������)
    // ============================================================

    // �����㹻����ڴ����洢 hex �ļ�����
    reg     [11:0] ad_memory     [0:32767];
    integer        ad_index = 0;

    // ��λ�Ĵ�����16λ (2 Leading Zeros + 12 Data + 2 Trailing Zeros)
    reg     [15:0] spi_shift_reg;

    // ��ʼ������ȡ hex �ļ�
    initial begin
        // ע�⣺��ȷ�� ad_data.hex �ڷ������Ĺ���Ŀ¼��
        // ������汨���Ҳ����ļ����볢��ʹ�þ���·�������� "D:/FPGA_Project/ad_data.hex"
        $readmemh("E:/pythonProject1/ad_data.hex", ad_memory);
        ad_in = 1'b0;
    end

    // ״̬������ CS �½��ؼ�����һ������x
    // �������߼�����ϵͳ�����������壨T0��ʱ��ǿ�Ƹ�λ��ȡ����
    always @(posedge u_dut.inst4_Order_4s.sys_start_pulse) begin
        ad_index = 0;
        $display("[%0t] AD Simulation Model: Reset ad_index to 0 (New Cycle Start)", $time);
    end


    // �������߼����� CS �½��أ����俪ʼ�����ص�ǰ���������ݵ���λ�Ĵ���
    always @(negedge ad_cs) begin
        // ���� 16 λ����֡��2λǰ��0 + 12λ���� + 2λ��׺0
        // AD7352 ��Ҫ 16 ��ʱ�����ڣ�����λ���м�
        if (ad_index < 32768) begin
            // ����ĸ�ʽ {2'b00, data, 2'b00} ��Ӧ AD.v �еĽ����߼�
            spi_shift_reg <= {2'b00, ad_memory[ad_index], 2'b00};

            // ׼����һ�ζ�ȡ������
            ad_index <= ad_index + 1;
        end
        else begin
            spi_shift_reg <= 16'd0;  // ���ݶ������ 0
        end

        $display("[%0t] AD Model: Loaded Data[%0d] = %h", $time, ad_index, ad_memory[ad_index]);
    end


    // ������λ��� (SPI Slave)
    // AD7352 �� SCLK �½��ظı����ݣ�FPGA (Master) �� SCLK �����ز���
    // ����� ad_clk �� FPGA �� AD.v ����
    always @(negedge ad_clk) begin
        if (!ad_cs) begin
            // ������λ
            ad_in <= spi_shift_reg[15];
            // ����
            spi_shift_reg <= {spi_shift_reg[14:0], 1'b0};
        end
        else begin
            ad_in <= 1'b0;
        end
    end

    // ============================================================
    // 9. ����������
    // ============================================================
    initial begin
        // --- ��ʼ�� ---
        rst_n = 1;
        TBS_in = 1;
        ad_index = 0;

        // --- ��λ & �ȴ� PLL �ȶ� ---
        #200;
        rst_n = 0;
        #200;
        rst_n = 1;
        #1000;

        $display("==================================================");
        $display("Simulation Start: Ultrasound System");
        $display("Data Source: ad_data.hex");
        $display("Simulating 10ms cycle...");
        $display("==================================================");

        // ========================================================
        // �׶� 1: ������������ 0x01
        // ========================================================
        $display("[%0t] Sending Command 0x01 (System Start)...", $time);
        send_tbs_byte(8'h01);

        // �ȴ�����������
        wait (debug_command == 3'h1);
        $display("[%0t] Command Received. System Starting...", $time);

        // ========================================================
        // �׶� 2: ���� 10ms ����
        // ========================================================
        // ��ʱ Order_4s ���� SYS_START -> WAIT_10MS
        // ������ PULSE_GEN (���䳬����) -> WAIT_1MS -> AD_SAMPLING
        // �� AD_SAMPLING �׶Σ�ad_cs ���᲻�Ϸ�ת����ȡ ad_data.hex �е�����

        // ���������㹻����ʱ�� (12ms) �Ը������� 10ms ���ڼ���������
        #12_000_000;

        // $display("==================================================");
        // $display("[%0t] Simulation Finished.", $time);
        // $display("Please check waveform for 'ad_in', 'ad_cs' and 'debug_ad_out_data'.");
        // $display("==================================================");
        // $stop;
    end

endmodule
