`timescale 1ns / 1ps // �������ʱ�䵥λΪ1ns������Ϊ1ps [1]
module tb_TBS_RX; // Testbench ģ��û����������˿� [1]
    // -- �������� --
    localparam CLK_FREQ    = 50_000_000;   // ʱ��Ƶ�� 50MHz
    localparam BAUD_RATE   = 115200;       // ������ 115200
    localparam CLK_PERIOD  = 1_000_000_000 / CLK_FREQ; // ʱ������: 20ns
    localparam BIT_PERIOD  = 1_000_000_000 / BAUD_RATE; // ��������: ~8680ns
    localparam PULSE_WIDTH = BIT_PERIOD / 10;          // TBS '0' ������: ~868ns
    // -- �źŶ��� --
    // DUT �����ź�����Ϊ reg
    reg clk_50M;
    reg rst_n;
    reg TBS_in;
    // DUT ����ź�����Ϊ wire
    wire rs232_out;
    
    //----------------------------------------------------------------
    // ��������ģ�� (DUT: Design Under Test)
    //----------------------------------------------------------------
    TBS_RX #(
        .CLK_FREQ(CLK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) u_tbs_rx (
        .clk_50M(clk_50M),
        .rst_n(rst_n),
        .TBS_in(TBS_in),
        .rs232_out(rs232_out)
    );
    //----------------------------------------------------------------
    // 1. ʱ�Ӻ͸�λ��������
    //----------------------------------------------------------------
    // ����ʱ���ź�
    initial begin
        clk_50M = 0;
        forever #(CLK_PERIOD / 2) clk_50M = ~clk_50M; // ��������Ϊ CLK_PERIOD ��ʱ��
    end
    // ���ɸ�λ�źźͲ���������
    initial begin
        // ��ʼ���͸�λ
        rst_n = 1'b0; // ���븴λ״̬
        TBS_in = 1'b1; // ���߿���Ϊ��
        #200;          // ���ָ�λ 200ns [3]
        rst_n = 1'b1; // �ͷŸ�λ
        #200;          // �ȴ���·�ȶ�
        $display("------------------- Simulation Start -------------------");
        
        // �������񣬷��Ͳ�������
        send_tbs_byte(8'h55); // ���� 01010101
        send_tbs_byte(8'hA3); // ���� 10100011
        send_tbs_byte(8'h00); // ����ȫ 0
        send_tbs_byte(8'hFF); // ����ȫ 1
        
        #50000; // �ȴ����һ���ֽڷ������
        
        $display("------------------- Simulation_Finish -------------------");
        $finish; // ��������
    end
    //----------------------------------------------------------------
    // 2. ������������ (Stimulus)
    //----------------------------------------------------------------
    // ����һ���������ڷ���һ���ֽڵ� TBS ��ʽ����
    task send_tbs_byte;
        input [7:0] data_to_send;
        integer i;
        begin
            $display("At time %0t ns, sending TBS byte: 0x%h", $time, data_to_send);
            
            // -- ������ʼλ (ֵΪ'0') --
            TBS_in = 1'b0;
            #(PULSE_WIDTH);
            TBS_in = 1'b1;
            #(BIT_PERIOD - PULSE_WIDTH);
            // -- ����8λ����λ (�ӵ�λ����λ) --
            for (i = 0; i < 8; i = i + 1) begin
                if (data_to_send[i] == 1'b0) begin
                    // ����� '0', ����һ��������
                    TBS_in = 1'b0;
                    #(PULSE_WIDTH);
                    TBS_in = 1'b1;
                    #(BIT_PERIOD - PULSE_WIDTH);
                end else begin
                    // ����� '1', ���ָߵ�ƽ
                    TBS_in = 1'b1;
                    #(BIT_PERIOD);
                end
            end
            // -- ����ֹͣλ (ֵΪ'1') --
            TBS_in = 1'b1;
            #(BIT_PERIOD);
            
            // �����ֽ�֮������һЩ����ʱ��
            #(BIT_PERIOD * 2);
        end
    endtask
    //----------------------------------------------------------------
    // 3. ��غͱȽ� (Monitor)
    //----------------------------------------------------------------
    // ��عؼ��źţ����źű仯ʱ��ӡ��״̬
    initial begin
        // $time �����ڻ�ȡ��ǰ����ʱ�� [1]
        $monitor("At time %0t ns: rst_n=%b, TBS_in=%b ===> rs232_out=%b",
                 $time, rst_n, TBS_in, rs232_out);
    end
endmodule
