`timescale 1ns / 1ps

module tb_Order_4s();

    // �����ź�
    reg        clk_50M;
    reg        rst_n;
    reg [2:0]  command;

    // ����ź�
    wire       start;
    wire       start_test;
    wire       Exc_start;
    wire       AD_start;

    // ʵ��������ģ��
    Order_4s uut (
        .clk_50M(clk_50M),
        .rst_n(rst_n),
        .command(command),
        .start(start),
        .start_test(start_test),
        .Exc_start(Exc_start),
        .AD_start(AD_start)
    );

    // ���� 50MHz ʱ��
    always #10 clk_50M = ~clk_50M;  // ���� 20ns �� 50MHz

    // ��ʼ��
    initial begin
        // ��ʼ���ź�
        clk_50M = 0;
        rst_n = 0;
        command = 3'h0;

        // �ͷŸ�λ
        #100;
        rst_n = 1;

        // ������������
        #50;
        command = 3'h1;  // ϵͳ����
        #50;
        command = 3'h0;  // �����źŽ���

        // ���� 1 ��
        #1000000000;  // 1 �� = 1,000,000,000 ns

        // ��������
        $display("Simulation finished at 1 second.");
        $finish;
    end

    // // ����źű仯
    // initial begin
    //     $monitor("Time = %t ns | State = %d | Command = %h | Start = %b | Exc_start = %b | AD_start = %b",
    //              $time, uut.current_state, command, start, Exc_start, AD_start);
    // end

    // ���� VCD �ļ����ڲ��η���
    initial begin
        $dumpfile("Order_4s.vcd");
        $dumpvars(0, tb_Order_4s);
    end

endmodule
