// `timescale 1ns / 1ps

// module tb_90khz;

//     // Parameters
//     parameter CLK_PERIOD = 20; // 50MHz clock period (20ns)
//     parameter SIM_TIME = 1_000_000_000; // 1 second simulation time

//     // Inputs
//     reg clk_50M;
//     reg rst_n;

//     // Outputs
//     wire VIN_1;
//     wire VIN_2;
//     wire VIN_3;
//     wire VIN_4;

//     // Instantiate the module
//     ultrasound_launch_90KHz_10ms uut (
//         .clk_50M(clk_50M),
//         .rst_n(rst_n),
//         .VIN_1(VIN_1),
//         .VIN_2(VIN_2),
//         .VIN_3(VIN_3),
//         .VIN_4(VIN_4)
//     );

//     // Clock generation
//     initial begin
//         clk_50M = 0;
//         forever #(CLK_PERIOD/2) clk_50M = ~clk_50M;
//     end

//     // Test sequence
//     initial begin
//         // Initialize signals
//         rst_n = 0;

//         // Reset the system
//         #(CLK_PERIOD*10) rst_n = 1; // Release reset after 10 clock cycles
//         #(CLK_PERIOD*10) rst_n = 0; // Assert reset again for a short duration
//         #(CLK_PERIOD*10) rst_n = 1; // Release reset

//         // Run the simulation for 1 second
//         #(SIM_TIME) $stop; // Stop simulation after 1 second
//     end

// endmodule
`timescale 1ns/1ps

module tb_90khz;

    // ʱ�Ӻ͸�λ�ź�
    reg clk_50M;
    reg rst_n;
    reg launch_cmd;
    
    // ����ź�
    wire VIN_1;
    wire VIN_2;
    wire VIN_3;
    wire VIN_4;
    
    // ʱ�Ӳ���
    parameter CLK_PERIOD = 20; // 50MHzʱ�ӣ�����20ns
    
    // ʵ����������ģ��
    ultrasound_launch_90KHz_10ms uut (
        .clk_50M(clk_50M),
        .rst_n(rst_n),
        .launch_cmd(launch_cmd),
        .VIN_1(VIN_1),
        .VIN_2(VIN_2),
        .VIN_3(VIN_3),
        .VIN_4(VIN_4)
    );
    
    // ʱ������
    always #(CLK_PERIOD/2) clk_50M = ~clk_50M;
    
    // ��ʼ��
    initial begin
        // ��ʼ���ź�
        clk_50M = 0;
        rst_n = 0;
        launch_cmd = 0;
        
        
        // ��λ����
        #100;
        rst_n = 1;
        #100;
        
        $display("=== ����������ģ����濪ʼ ===");
        $display("ʱ��: %t", $time);
        
        // ���Գ���1�����η���
        $display("\n--- ����1�����η��� ---");
        launch_cmd = 1;
        #20; // �ȴ�20ns
        launch_cmd = 0;
        #10000000; // �ȴ�10ms
        
        // ���Գ���2���������ٷ��䣨ģ������������
        $display("\n--- ����2���������� ---");
        repeat (3) begin
            launch_cmd = 1;
            #200000; // 200us
            launch_cmd = 0;
            #5000000; // 5ms���
        end
        
        // ���Գ���3����ʱ�䱣�ַ���
        $display("\n--- ����3����ʱ�䷢�� ---");
        launch_cmd = 1;
        #5000000; // 5ms
        launch_cmd = 0;
        #10000000; // 10ms
        
        // ���Գ���4����λ����
        $display("\n--- ����4����λ���� ---");
        rst_n = 0;
        #1000;
        rst_n = 1;
        #1000000;
        
        // ���Գ���5���߽��������
        $display("\n--- ����5���߽�������� ---");
        launch_cmd = 1;
        #100;
        launch_cmd = 0;
        #100000;
        launch_cmd = 1;
        #1000000;
        launch_cmd = 0;
        
        // �ȴ�ʣ��ʱ�����100ms����
        #80000000; // 80ms
        
        $display("\n=== ������� ===");
        $display("�ܷ���ʱ��: %t", $time);
        $finish;
    end
    
    // �������ź�
    integer vin1_count = 0;
    integer vin2_count = 0;
    integer vin3_count = 0;
    integer vin4_count = 0;
    reg vin1_last = 0;
    reg vin2_last = 0;
    reg vin3_last = 0;
    reg vin4_last = 0;
    
    always @(posedge clk_50M) begin
        // ͳ��VIN_1��������
        if (VIN_1 && !vin1_last) begin
            vin1_count <= vin1_count + 1;
        end
        vin1_last <= VIN_1;
        
        // ͳ��VIN_2��������
        if (VIN_2 && !vin2_last) begin
            vin2_count <= vin2_count + 1;
        end
        vin2_last <= VIN_2;
        
        // ͳ��VIN_3��������
        if (VIN_3 && !vin3_last) begin
            vin3_count <= vin3_count + 1;
        end
        vin3_last <= VIN_3;
        
        // ͳ��VIN_4��������
        if (VIN_4 && !vin4_last) begin
            vin4_count <= vin4_count + 1;
        end
        vin4_last <= VIN_4;
    end
    
    

endmodule
