`timescale 1ns/1ns

module tb_Echo;

    // ============================================================
    // 1. ��������
    // ============================================================
    parameter CLK_PERIOD = 20;      // 50MHzʱ������ = 20ns
    parameter AD_SAMPLE_RATE = 50;  // 1MHz������ = 50��ʱ������
    parameter DATA_DEPTH = 5000;    // �����������

    // ============================================================
    // 2. �źŶ���
    // ============================================================
    reg clk_50M;
    reg rst_n;
    
    // ����������Ӧ Echo.vhd �Ķ�������
    reg sys_start_pulse;    // ��ע�⡿��Ҫ�� BDF/VHDL �в�������˿�
    reg [17:0] corr_threshold; // ��ע�⡿��Ҫ�� BDF/VHDL �в�������˿�
    
    reg ad_valid_in;        // ��Ӧ DSP ������ valid
    reg [11:0] ad_data_in;  // ��Ӧ DSP ������ data (ԭʼ12λ)

    // ����ź�
    wire [31:0] echo_tof;
    wire [17:0] echo_peak;
    wire hit_flag;
    wire signed [12:0] debug_clean_data; 
    wire signed [31:0] debug_dsp_sum;    // �鿴 DSP �ڲ��ۼ�����ԭʼֵ
    
    assign debug_clean_data = uut.dsp_data_wire; 
    assign debug_dsp_sum    = uut.u_dsp.sum;     // ��������ֱ�ӿ���ģ������źţ�
    // �洢�����飬���ڴ�� Hex ����
    reg [11:0] mem_data [0:DATA_DEPTH-1];
    integer i;

    // ============================================================
    // 3. ʵ��������ģ�� (Top Level: Echo)
    // ============================================================
    // ע�⣺������ VHDL ��û�м� start_pulse �� threshold������ᱨ��
    // ����ظ������ VHDL �ļ���
    Echo uut (
        .clk_50M(clk_50M), 
        .rst_n(rst_n), 
        
        // �ؼ������ź� (������ӵ�����)
        .sys_start_pulse(sys_start_pulse), 
        .corr_threshold(corr_threshold), 
        // ���������� (ι�� DSP)
        .ad_valid_in(ad_valid_in), 
        .ad_data_in(ad_data_in), 
        
        // ������
        .hit_flag(hit_flag), 
        .echo_peak(echo_peak), 
        .echo_tof(echo_tof)
    );

    // ============================================================
    // 4. ʱ������
    // ============================================================
    always #(CLK_PERIOD/2) clk_50M = ~clk_50M;

    // ============================================================
    // 5. �����Թ���
    // ============================================================
    initial begin
        // --- ��ʼ�� ---
        clk_50M = 0;
        rst_n = 0;
        sys_start_pulse = 0;
        ad_valid_in = 0;
        ad_data_in = 0;
        
        // ������ֵ�����ھ��� FIR �˲����źŷ�ֵ���ܱ仯��
        // ���������һ��۲죬���߸��� DSP �ڲ��ضϺ�Ĳ��ε���
        corr_threshold = 18'd1000; 

        // --- ���������ļ� ---
        // ·�������ʵ������޸�
        $readmemh("E:/pythonProject1/ad_data.hex", mem_data);
        $display("Data loaded from ad_data.hex");

        // --- ��λ�ͷ� ---
        #100;
        rst_n = 1;
        #100;

        // --- ����ϵͳ�������� (T0ʱ��) ---
        @(posedge clk_50M);
        sys_start_pulse = 1;
        @(posedge clk_50M);
        sys_start_pulse = 0;

        // --- ��ʼģ�� AD ������ (1MHz) ---
        // ע�⣺�������ǰ�����ι�� Echo ���� -> DSP -> Correlation
        for (i = 0; i < 4500; i = i + 1) begin
            // ģ�� AD ת������ź�
            @(posedge clk_50M);
            ad_valid_in = 1;
            ad_data_in = mem_data[i]; // ����ԭʼ 12λ ����
            
            @(posedge clk_50M);
            ad_valid_in = 0; 

            // �ȴ���һ��������
            repeat(AD_SAMPLE_RATE - 2) @(posedge clk_50M);

            // --- ʵʱ��ӡ������Ϣ ---
            // ע�⣺���� uut �� VHDL��uut.b2v_inst1 ���ڲ�ʵ��
            // ModelSim ��ͨ��֧�ֿ����Բ�����ã����������ע�͵������ display
            /* b2v_inst1 �� Echo.vhd ��ʵ������ echo_correlation ������
               sum/abs_sum �� echo_correlation �ڲ��ź�
               ����·�����ƿ�����Ҫ���� ModelSim �� Objects ����ȷ��
            */
             if (hit_flag) begin
                 $display("HIT! Time: %t | Index: %d | Peak: %d | ToF: %d", 
                          $time, i, echo_peak, echo_tof);
             end
        end

        // --- ������� ---
        #1000;
        $display("Simulation Finished.");
        $display("Final ToF: %d (x20ns)", echo_tof);
        $display("Final Peak: %d", echo_peak);
        $stop;
    end

endmodule