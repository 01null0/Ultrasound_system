`timescale 1ns/1ns

module tb_Echo_Correlation_SpeedTest;

    // ==========================================
    // 1. �������ò��� (�ڴ˴��޸��Բ��Բ�ͬ���)
    // ==========================================
    parameter CLK_PERIOD      = 20;     // 50MHz (20ns)
    parameter TEST_DATA_DEPTH = 5000;  // ���޸��������Ҫ���Ե������� (���� 2000, 10000, 50000)
    
    // Hex�ļ�·�� (�����ʵ������޸�)
    parameter HEX_FILE_PATH   = "E:/pythonProject1/ad_data.hex"; 

    // ==========================================
    // 2. �źŶ���
    // ==========================================
    reg clk_50M;
    reg rst_n;
    reg sys_start_pulse;

    // FIFO �ӿ�
    reg  [11:0] fifo_data_in;
    reg         fifo_wrreq;
    wire        fifo_rdreq;
    wire [11:0] fifo_q;
    wire        fifo_empty;
    
    // DUT ���
    reg  [17:0] corr_threshold;
    wire [19:0] echo_tof;
    wire [17:0] echo_peak;
    wire        hit_flag;
    wire        processing_done;

    // �洢�������
    reg [11:0] mem_data [0:100000]; // ȷ��������鹻����װ������Hex�ļ�
    integer i;
    
    // ��ʱͳ�Ʊ���
    time start_time;
    time end_time;
    integer process_cycles;

    // ==========================================
    // 3. ģ��ʵ����
    // ==========================================
    
    // 3.1 FIFO (ʹ���������е� FIFO)
    fifo u_fifo (
        .data    (fifo_data_in),
        .wrclk   (clk_50M),
        .wrreq   (fifo_wrreq),
        .rdclk   (clk_50M),
        .rdreq   (fifo_rdreq),
        .q       (fifo_q),
        .rdempty (fifo_empty)
    );

    // 3.2 ����ģ�� (DUT)
    Echo_Correlation uut (
        .clk_50M         (clk_50M), 
        .rst_n           (rst_n), 
        .sys_start_pulse (sys_start_pulse), 
        .fifo_q          (fifo_q),
        .fifo_empty      (fifo_empty),
        .fifo_rdreq      (fifo_rdreq),
        .corr_threshold  (corr_threshold), 
        .echo_tof        (echo_tof), 
        .echo_peak       (echo_peak), 
        .hit_flag        (hit_flag),
        .processing_done (processing_done)
    );

    // ==========================================
    // 4. ʱ������
    // ==========================================
    initial clk_50M = 0;
    always #(CLK_PERIOD/2) clk_50M = ~clk_50M;

    // ==========================================
    // 5. ���ܼ���߼� (��������)
    // ==========================================
    
    // ��ش���ʼ (�� FIFO ��һ�α���ȡʱ)
    reg measurement_started;
    initial measurement_started = 0;

    always @(posedge clk_50M) begin
        if (fifo_rdreq && !measurement_started) begin
            start_time = $time;
            measurement_started = 1;
            $display("[Time: %t] Processing STARTED.", $time);
        end
    end

    // ==========================================
    // 6. �����Լ��� (ȫ��д��)
    // ==========================================
    initial begin
        // --- ��ʼ�� ---
        rst_n = 0;
        sys_start_pulse = 0;
        fifo_wrreq = 0;
        fifo_data_in = 0;
        corr_threshold = 18'd2500; // ������ֵ
        
        // --- �������� ---
        // ע�⣺��ȷ�� Hex �ļ��е������� >= TEST_DATA_DEPTH
        $readmemh(HEX_FILE_PATH, mem_data);
        $display("--------------------------------------------------");
        $display("Test Configuration:");
        $display("  Data Depth: %d samples", TEST_DATA_DEPTH);
        $display("  Clock Freq: 50 MHz");
        $display("--------------------------------------------------");

        // --- ��λ�ͷ� ---
        #100;
        rst_n = 1;
        #100;
        
        // --- ���� Start Pulse (�����ڲ�������) ---
        @(posedge clk_50M);
        sys_start_pulse = 1;
        @(posedge clk_50M);
        sys_start_pulse = 0;
        
        // �ȴ���������
        repeat(5) @(posedge clk_50M);

        // --- ���ؼ���ȫ��д��ѭ�� ---
        $display("[Time: %t] Starting FAST WRITE to FIFO...", $time);
        
        for (i = 0; i < TEST_DATA_DEPTH; i = i + 2) begin 
            // ׼������
            fifo_data_in = mem_data[i]; // ����hex�ļ��������洢��
            fifo_wrreq = 1;
            
            // ÿ��ʱ������д��һ�����ݣ����ȴ���
            @(posedge clk_50M); 
        end
        
        // ֹͣд��
        fifo_wrreq = 0;
        fifo_data_in = 0;
        $display("[Time: %t] Fast Write COMPLETED. Waiting for DUT to finish...", $time);

        // --- �ȴ� FIFO ��ȡ�� ---
        // ֻҪ FIFO �ǿգ����� DUT ���������Ч��־��������ӳ٣����͵ȴ�
        // ����� fifo_empty ����ֱ�ӵ��о�
        wait(fifo_empty == 1);
        
        // �ٶ���ȴ�һС��ʱ�䣬ȷ����ˮ�����꣨���� 100�����ڣ�
        repeat(100) @(posedge clk_50M);
        
        end_time = $time;
        
        // --- ���ͳ�ƽ�� ---
        $display("--------------------------------------------------");
        $display("PERFORMANCE REPORT");
        $display("--------------------------------------------------");
        $display("Samples Processed : %d", TEST_DATA_DEPTH);
        $display("Total Time Taken  : %t ns", end_time - start_time);
        
        process_cycles = (end_time - start_time) / CLK_PERIOD;
        $display("Total Clock Cycles: %d", process_cycles);
        
        // ����ƽ���ٶ�
        // ���������Ӧ���� 1 cycle/sample
        $display("Average Speed     : %0.2f cycles/sample", (process_cycles * 1.0) / TEST_DATA_DEPTH);
        $display("--------------------------------------------------");

        if (hit_flag)
            $display("RESULT: Hit DETECTED at Index %d, Peak %d", echo_tof, echo_peak);
        else
            $display("RESULT: No Hit Detected.");

        $stop;
    end

endmodule
