module UART_RX (
    input             clk_50M,       // 50MHzʱ��
    input             rst_n,         // ��λ�ź�
    input             rs232_rx,      // ������������
    output reg        rx_done,       // ������ɱ�־
    output     [11:0] test_rx_data,  // ���յ�������
    output reg [ 2:0] command        // �������
);
    //��������
    parameter CLK_FREQ = 50_000_000;  // ϵͳʱ��Ƶ��
    parameter BAUD_RATE = 115200;  // ������
    //localparam BAUD_CNT_MAX = CLK_FREQ / BAUD_RATE - 1;  // �������ڼ��������ֵ
    //localparam HALF_BAUD = BAUD_CNT_MAX/2;  // �벨�����ڼ��㣨651��
    localparam BAUD_CNT_MAX = 434;
    localparam HALF_BAUD = 217;

    //�źŶ���
    reg [ 1:0] sync_regs;  // ͬ���Ĵ�������������̬������
    reg [16:0] baud_cnt;  // �����ʼ�����
    reg [ 3:0] bit_cnt;  // ����λ������
    reg        rx_en;  // ����ʹ���ź�
    reg [ 7:0] rx_data;
    assign test_rx_data = {4'b1010, rx_data};  //�������

    //״̬����
    localparam IDLE = 2'b00;  // ����״̬
    localparam START = 2'b01;  // ��ʼλ���
    localparam DATA = 2'b10;  // ����λ����
    localparam STOP = 2'b11;  // ֹͣλ����
    reg [1:0] state;

    //ͬ�����½��ؼ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) sync_regs <= 2'b11;
        else sync_regs <= {sync_regs[0], rs232_rx};
    end
    wire nedge_detect = (sync_regs[1] & ~sync_regs[0]);  // �½��ؼ��

    //��״̬��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            state    <= IDLE;
            baud_cnt <= 0;
            bit_cnt  <= 0;
            rx_data  <= 8'h00;
            rx_done  <= 0;
            rx_en    <= 0;
        end
        else begin
            if (rx_done) begin
                rx_done <= 1'b0;
                rx_data <= 0;
            end
            case (state)
                IDLE: begin
                    if (nedge_detect) begin  // ��⵽��ʼλ�½���
                        state <= START;
                        baud_cnt <= 0;
                    end
                end

                START: begin  // ��ʼλ��֤
                    if (baud_cnt == HALF_BAUD) begin  // �޸�ΪHALF_BAUD
                        if (!sync_regs[0]) begin  // ȷ����ʼλΪ��
                            state <= DATA;
                            baud_cnt <= 0;
                            bit_cnt <= 0;
                        end
                        else state <= IDLE;  // ���󣬷��ؿ���
                    end
                    else baud_cnt <= baud_cnt + 1;
                end

                DATA: begin  // ����8λ����
                    if (baud_cnt == BAUD_CNT_MAX) begin
                        baud_cnt <= 0;
                        if (bit_cnt == 7) begin
                            state <= STOP;
                        end
                        else bit_cnt <= bit_cnt + 1;
                    end
                    else begin
                        if (baud_cnt == HALF_BAUD) begin  // �޸�ΪHALF_BAUD
                            rx_data[bit_cnt] <= sync_regs[0];  // �ڱ����м����
                        end
                        baud_cnt <= baud_cnt + 1;
                    end
                end

                STOP: begin  // ֹͣλ����
                    if (baud_cnt == BAUD_CNT_MAX) begin
                        if (sync_regs[0] == 1'b1) begin  // ��ֹ֤ͣλΪ��
                            rx_done <= 1'b1;  // ���ݽ������
                        end
                        state <= IDLE;
                    end
                    else baud_cnt <= baud_cnt + 1;
                end
            endcase
        end
    end

    //�������
    wire [7:0] cmd = rx_data;
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            command <= 0;
        end
        else begin
            if (rx_done) begin
                case (cmd)
                    8'h00: command <= 0;
                    8'h01: command <= 1;
                    8'h02: command <= 2;
                    8'h03: command <= 3;
                    8'h04: command <= 4;
                    8'h05: command <= 5;
                    8'h06: command <= 6;
                    8'h07: command <= 7;
                    8'h08: command <= 8;

                    default: command <= 0;
                endcase
            end
            else begin

                command <= 0;
            end
        end
    end
endmodule
