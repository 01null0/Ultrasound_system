// ϵͳ������ʼ4���ʱ
// ÿ10ms����һ�γ�������
// �������ӳ�1ms��ʼAD����
// AD��������8ms��1ms-9ms�ڼ䣩
// 4���ϵͳ�Զ�ֹͣ
module Order (
    input            clk_50M,     // 50MHzʱ��
    input            rst_n,       // ��λ�ź�
    input      [2:0] command,     // ��������
    output reg       start,       // ϵͳ����
    output reg       start_test,  // ��ʼ����
    output reg       Exc_start,   //������ʼ�ź�
    output reg       AD_start     //AD��ʼ�ź�
    // ,output reg       AD_end       //ADֹͣ�źţ���ʱҲ����ϵͳֹͣ
);
    //��������
    parameter CLK_FREQ = 50_000_000;  // ϵͳʱ��Ƶ��
    parameter Time_4s = 200_000_000;  // 4S
    parameter Time_10ms = 500_000;  // 10mS
    parameter Time_9ms = 450_000;  // 9ms
    parameter Time_1ms = 50_000;  // 1ms
    parameter Time_1us = 50;  // 4S

    reg [27:0] cnt_4s;  //4s������
    reg [18:0] cnt_10ms;  //10ms������
    reg [ 5:0] cnt_1us;  //1us������
    reg        cnt_en;  //4s����ʱ���ź�ʹ��
    reg [ 1:0] sync_regs;  // ͬ���Ĵ�������������̬������
    reg [ 1:0] sync_regs_test;
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            start <= 0;
            start_test <= 0;
        end
        else begin
            case (command)
                3'h0: begin
                    start <= 0;
                    start_test <= 0;
                end
                3'h1: start <= 1;  //ϵͳ������������ʱ��
                3'h2: start_test <= 1;  //����������������ʱ��
                default: begin
                    start <= 0;
                    start_test <= 0;
                end
            endcase
        end
    end

    //ͬ�����½��ؼ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) sync_regs <= 2'b11;
        else sync_regs <= {sync_regs[0], start};
    end
    wire nedge_detect = (sync_regs[1] & ~sync_regs[0]);  // �����ź�start�½��ؼ��

    //ͬ�����½��ؼ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) sync_regs_test <= 2'b11;
        else sync_regs_test <= {sync_regs_test[0], start_test};
    end
    wire nedge_detect_test = (sync_regs_test[1] & ~sync_regs_test[0]);  // �����ź�start_test�½��ؼ��

    //�����趨4S��Ϊ�ɼ�ʱ�䣬���ಿ��Ϊ�����������ʱ������

    //4s��ʱ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            cnt_4s <= Time_4s + 1;
            cnt_en <= 0;
        end
        else if (cnt_4s == Time_4s) begin
            cnt_4s <= Time_4s + 1;
            cnt_en <= 0;
        end
        else if (nedge_detect) begin
            cnt_4s <= 0;
        end
        else begin
            cnt_4s <= cnt_4s + 1;
            cnt_en <= 1;
        end
    end
    //10ms��ʱ�������ڼ��������ź�
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            cnt_10ms <= Time_10ms + 1;
        end
        else if (!cnt_en) begin
            cnt_10ms <= Time_10ms + 1;
        end
        else if (cnt_10ms == Time_10ms) begin
            cnt_10ms <= 0;
        end
        else if (nedge_detect) begin
            cnt_10ms <= 0;
        end
        else begin
            cnt_10ms <= cnt_10ms + 1;
        end
    end

    //90KHZ��ʮ�������ʣ����ô���1MHZ������
    //1us��ʱ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            cnt_1us <= Time_1us + 1;
        end
        else if (!cnt_en) begin
            cnt_1us <= Time_1us + 1;
        end
        else if (cnt_1us == Time_1us) begin
            cnt_1us <= 0;
        end
        else if (cnt_10ms == Time_1ms) begin
            cnt_1us <= 0;  //�������1ms�󣬿���ADת��
        end
        else if (cnt_10ms == Time_9ms) begin
            cnt_1us <= Time_1us + 1;
        end
        else begin
            cnt_1us <= cnt_1us + 1;
        end
    end

    //4s�����󣬷���ֹͣ�ź�
    // always @(posedge clk_50M or negedge rst_n) begin
    //     if (!rst_n) begin
    //         AD_end <= 0;
    //     end
    //     else if (cnt_4s == Time_4s) begin
    //         AD_end <= 1;
    //     end
    //     else begin
    //         AD_end <= 0;
    //     end
    // end

    //10ms����һ�γ�������
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            Exc_start <= 0;
        end
        else if (cnt_10ms == Time_10ms) begin
            Exc_start <= 1;
        end
        else begin
            Exc_start <= 0;
        end
    end
    //������ɺ�1ms��ʼAD�ɼ�
    //ÿ��1us��AD����һ��
    always @(posedge clk_50M or negedge rst_n) begin
        if (!rst_n) begin
            AD_start <= 0;
        end
        else if (cnt_1us == Time_1us) begin
            AD_start <= 1;
        end
        else begin
            AD_start <= 0;
        end
    end

endmodule
