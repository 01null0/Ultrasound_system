`timescale 1ns / 1ps

module tb_UART_RX();
    // �����ź�
    reg clk_50M;
    reg rst_n;
    reg rs232_rx;
    
    // ����ź�
    wire rx_done;
    //wire [7:0] rx_data;
    wire [2:0] command;
    parameter BPS=8681;// 1/38400�� �� 26041ns
    // ʵ����UART_RXģ��
    UART_RX uut (
        .clk_50M(clk_50M),
        .rst_n(rst_n),
        .rs232_rx(rs232_rx),
        .rx_done(rx_done),
        //.rx_data(rx_data),
        .command(command)
    );
    
    // ʱ�����ɣ�50MHz
    always #10 clk_50M = ~clk_50M;
    
    // ���񣺷���һ���ֽ�
    task send_byte;
        input [7:0] data;
        integer i;
        begin
            // ��ʼλ
            rs232_rx = 0;
            #BPS; 
            
            // ����λ
            for (i = 0; i < 8; i = i + 1) begin
                rs232_rx = data[i];
                #BPS;
            end
            
            // ֹͣλ
            rs232_rx = 1;
            #BPS;
        end
    endtask
    
    // ��������
    initial begin
        // ��ʼ���ź�
        clk_50M = 0;
        rst_n = 0;
        rs232_rx = 1; // ����״̬Ϊ�ߵ�ƽ
        
        // ��λ
        #100 rst_n = 1;
        
        // �ȴ�һ��ʱ��
        #1000;
        
        // ����1����������0x01
        send_byte(8'h01);
        
        // �ȴ��������
        #100000;
        
        // ����2����������0x02
        send_byte(8'h02);
        
        // �ȴ��������
        #100000;
        
        // ����3����������0x04
        send_byte(8'h04);
        
        // �ȴ��������
        #100000;
        
        // ����4��������Ч����
        send_byte(8'hFF);
        
        // �ȴ��������
        #100000;
        
        // ��������
        #100 $finish;
    end
    
endmodule
