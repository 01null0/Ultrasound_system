`timescale 1ns/1ns

module tb_Echo_Correlation;

    // ==========================================
    // 1. ��������
    // ==========================================
    parameter CLK_PERIOD = 20;      // 50MHzϵͳʱ�� (20ns)
    // ģ�� ADC �����ʣ�����Ϊ 1MHz (ÿ50��ϵͳʱ��дһ��FIFO)
    // �����Ը���ʵ���������д���ٶȣ��ⲻ��Ӱ�촦��������Ϊ�����ǻ�������������
    parameter ADC_WRITE_DELAY = 50; 
    
    parameter DATA_DEPTH = 20000;   // �����������

    // ==========================================
    // 2. �źŶ���
    // ==========================================
    reg clk_50M;
    reg rst_n;
    reg sys_start_pulse;
    
    // --- FIFO ����ź� ---
    reg  [11:0] fifo_data_in;   // д��FIFO������ (ģ��ADC���)
    reg         fifo_wrreq;     // FIFOд����
    wire        fifo_rdreq;     // FIFO������ (����DUT)
    wire [11:0] fifo_q;         // FIFO�������� (�͸�DUT)
    wire        fifo_empty;     // FIFO�ձ�־
    // -------------------

    // --- DUT ��������� ---
    reg  [17:0] corr_threshold;
    wire [19:0] echo_tof;       // �������������
    wire [17:0] echo_peak;
    wire        hit_flag;
    wire        processing_done; // ָʾFIFO�������

    // �洢������ (Hex�ļ�����)
    reg [11:0] mem_data [0:DATA_DEPTH-1];
    integer i;

    // ==========================================
    // 3. ģ��ʵ����
    // ==========================================

    // (1) ʵ���� FIFO (ʹ���������е� project/FIFO/fifo.v)
    // ע�⣺����ʱ��Ҫ���� fifo.v ���������� Altera ��
    fifo u_fifo (
        .data    (fifo_data_in),
        .wrclk   (clk_50M),      // ģ��дʱ��
        .wrreq   (fifo_wrreq),
        
        .rdclk   (clk_50M),      // ϵͳ��ʱ��
        .rdreq   (fifo_rdreq),
        .q       (fifo_q),
        .rdempty (fifo_empty)
    );

    // (2) ʵ��������ģ�� (Echo_Correlation_FIFO)
    Echo_Correlation uut (
        .clk_50M         (clk_50M), 
        .rst_n           (rst_n), 
        .sys_start_pulse (sys_start_pulse), 
        
        // FIFO �ӿ�����
        .fifo_q          (fifo_q),
        .fifo_empty      (fifo_empty),
        .fifo_rdreq      (fifo_rdreq),
        
        .corr_threshold  (corr_threshold), 
        .echo_tof        (echo_tof), 
        .echo_peak       (echo_peak), 
        .hit_flag        (hit_flag),
        .processing_done (processing_done)
    );

    // ==========================================
    // 4. ʱ������
    // ==========================================
    initial clk_50M = 0;
    always #(CLK_PERIOD/2) clk_50M = ~clk_50M;

    // ==========================================
    // 5. �����Լ���
    // ==========================================
    initial begin
        // --- ��ʼ�� ---
        rst_n = 0;
        sys_start_pulse = 0;
        fifo_wrreq = 0;
        fifo_data_in = 0;
        
        // ������ֵ (��������Hex���ݵ���)
        corr_threshold = 18'd4500; 

        // --- �������� ---
        // ������ԭ���� hex �ļ�·������
        $readmemh("E:/pythonProject1/ad_data.hex", mem_data);
        $display("Data loaded from ad_data.hex");

        // --- ��λ�ͷ� ---
        #100;
        rst_n = 1;
        #100;

        // --- ����ϵͳ�������� ---
        // �������ģ���ڵķ�ֵ��¼�ͼ�����
        @(posedge clk_50M);
        sys_start_pulse = 1;
        @(posedge clk_50M);
        sys_start_pulse = 0;

        $display("Starting to fill FIFO...");

        // --- ģ�� ADC ����д�� FIFO ---
        // ѭ����ȡ mem_data ��д�� FIFO
        for (i = 0; i < DATA_DEPTH; i = i + 1) begin // ע�⣺��������� +1 �� +2��ȡ�����������ݴ洢��ʽ
            
            // 1. ׼������
            fifo_data_in = mem_data[i];
            
            // 2. ����д��������
            @(posedge clk_50M);
            fifo_wrreq = 1;
            
            @(posedge clk_50M);
            fifo_wrreq = 0; // дʹ������
            
            // 3. ģ��������
            // ���� 1MHz �����ʣ�����Ҫ�ȴ�Լ 50 ��ʱ��������д��һ��
            // �������ģ�⡰�ȴ洢�����������������ʱ�ǳ�С�����ٰ�FIFO����
            repeat(ADC_WRITE_DELAY - 1) @(posedge clk_50M);
            
            // (��ѡ) ��ӡ����
            if (i % 1000 == 0) $display("Written sample %d to FIFO", i);
        end

        $display("All data written to FIFO.");
        
        // �ȴ� FIFO ��������
        wait(fifo_empty == 1);
        #1000; // �ٶ��һ���ȷ�����Ĵ������
        
        $stop;
    end

    // ==========================================
    // 6. ������ (��ѡ)
    // ==========================================
    // always @(posedge clk_50M) begin
    //     if (hit_flag) begin
    //         $display("Hit Detected! Sample Index: %d, Peak: %d", echo_tof, echo_peak);
    //     end
    // end

endmodule
