module FIFO_Buffer (
    input         clk,          // 50MHz
    input         rst_n,
    
    // д�ӿ� (���� AD)
    input         wr_en,        // AD ����ź� (ad_done)
    input  [11:0] wr_data,      // AD ���� (ad_out)
    output        full,         // �������ˣ�֪ͨ Order_4s ֹͣ����
    
    // ���ӿ� (���� UART)
    input         rd_req,       // UART ����ʱ�����ȡ
    output [11:0] rd_data,      // ���͸� UART ������
    output reg    rd_valid,     // ����������Ч (��Ϊ UART �� ad_done)
    output        empty         // �������
);

    // ���建����ȣ�4096 ���� (ռ�� EP4CE10 Լ 12% ���ڴ�)
    parameter DEPTH = 4096;
    parameter ADDR_W = 12; // 2^12 = 4096

    reg [11:0] mem [0:DEPTH-1]; // ���� RAM
    reg [ADDR_W-1:0] wr_ptr;
    reg [ADDR_W-1:0] rd_ptr;
    reg [ADDR_W:0]   cnt;       // ������������

    assign full  = (cnt >= DEPTH);
    assign empty = (cnt == 0);
    assign rd_data = mem[rd_ptr]; // ��������

    // д�߼�
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            wr_ptr <= 0;
        end else if (wr_en && !full) begin
            mem[wr_ptr] <= wr_data;
            wr_ptr <= wr_ptr + 1;
        end
    end

    // ���߼�
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rd_ptr <= 0;
            rd_valid <= 0;
        end else begin
            rd_valid <= 0; // Ĭ������
            if (rd_req && !empty) begin
                rd_ptr <= rd_ptr + 1;
                rd_valid <= 1; // ����һ��������� UART ���ݺ���
            end
        end
    end

    // �������߼�
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cnt <= 0;
        end else begin
            case ({wr_en && !full, rd_req && !empty})
                2'b10: cnt <= cnt + 1; // ֻд
                2'b01: cnt <= cnt - 1; // ֻ��
                default: cnt <= cnt;   // ͬʱ��д���޲���
            endcase
        end
    end

endmodule
